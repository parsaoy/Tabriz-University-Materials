module FourBitFullAdder(input [3:0]X,input[3:0]Y ,output [4:0] s);

	assign s=X+Y;

endmodule
library verilog;
use verilog.vl_types.all;
entity Comparator is
end Comparator;

library verilog;
use verilog.vl_types.all;
entity tbMemory is
end tbMemory;

library verilog;
use verilog.vl_types.all;
entity tbPriority_Encoder83 is
end tbPriority_Encoder83;

module SampleVerilog(X,Y);
	input X;
	output Y;
	not not1(Y,X);

endmodule
library verilog;
use verilog.vl_types.all;
entity tbDecoder24_DataFlow is
end tbDecoder24_DataFlow;

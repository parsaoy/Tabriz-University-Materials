library verilog;
use verilog.vl_types.all;
entity tbDecoder24_GateLevel is
end tbDecoder24_GateLevel;

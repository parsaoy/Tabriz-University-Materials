module adjoints(input [2:0] A, input B, output F);

if({A,B} == 4'b0011)
	{F = 1
	}
endmodule
library verilog;
use verilog.vl_types.all;
entity Display_Monitor is
end Display_Monitor;

module subtractModule(input [3:0]X, input [3:0]Y,output [4:0] T);

	assign T = X-Y;
	
endmodule
library verilog;
use verilog.vl_types.all;
entity tbBinaryToCommonAnode7Seg is
end tbBinaryToCommonAnode7Seg;

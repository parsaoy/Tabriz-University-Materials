library verilog;
use verilog.vl_types.all;
entity tbEightBitShiftRegiter is
end tbEightBitShiftRegiter;
